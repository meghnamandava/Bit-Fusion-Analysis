module fixed4 #(parameter COL_WIDTH=11) (
    input [7:0] in,
    input [7:0] weight,
    input [(COL_WIDTH*2)-1:0] psum_in,
    input s_in,
    input s_weight,
    output reg [(COL_WIDTH*2)-1:0] psum_fwd
    );

    always @(*) begin
        if (s_in == 1'b1 && s_weight == 1'b1) begin
            psum_fwd <= $signed(in[3:0]) * $signed(weight[3:0]) + $signed(in[7:4]) * $signed(weight[7:4]) + psum_in
        end else if (s_in == 1'b1 && s_weight == 1'b0) begin
            psum_fwd <= ($signed(in[3:0]) * weight[3:0]) + ($signed(in[7:4]) * weight[7:4]) + psum_in;
        end else if (s_in == 1'b0 && s_weight == 1'b1) begin
            psum_fwd <= (in[3:0] * $signed(weight[3:0])) + (in[7:4] * $signed(weight[7:4])) + psum_in;
        end else if (s_in == 1'b0 && s_weight== 1'b0) begin
            psum_fwd <= (in[3:0] * weight[3:0]) + (in[7:4] * weight[7:4]) + psum_in;
        end
    end    

 
endmodule

    