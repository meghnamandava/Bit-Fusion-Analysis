`timescale 1ns/1ns

module accelerator #(parameter ARRAY_SIZE=8) 
    (

    input clk, 
    input rst);

endmodule    